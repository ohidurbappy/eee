* C:\Users\Bappy\Desktop\PSpiceSchematics\Schematic4.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 25 11:00:00 2018



** Analysis setup **
.DC LIN V_V1 .5 20 1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic4.net"
.INC "Schematic4.als"


.probe


.END
