* C:\Users\Bappy\Desktop\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Tue Jul 17 08:58:54 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
