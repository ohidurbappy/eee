* C:\Users\Bappy\Desktop\PSpiceSchematics\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 25 10:25:59 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
