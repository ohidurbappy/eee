* C:\Users\Bappy\Desktop\Schematic5.sch

* Schematics Version 9.1 - Web Update 1
* Tue Jul 17 10:05:18 2018



** Analysis setup **
.DC LIN V_V1 1V 10V 2 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic5.net"
.INC "Schematic5.als"


.probe


.END
