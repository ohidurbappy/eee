* C:\Users\Bappy\Desktop\Schematic\Schematic8.sch

* Schematics Version 9.1 - Web Update 1
* Tue Jul 24 11:34:25 2018



** Analysis setup **
.DC LIN V_V1 0 20 2 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic8.net"
.INC "Schematic8.als"


.probe


.END
