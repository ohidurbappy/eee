* C:\Users\Bappy\Desktop\PSpiceSchematics\Schematic10.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 25 11:54:22 2018



** Analysis setup **
.tran 0ns 0.1s
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic10.net"
.INC "Schematic10.als"


.probe


.END
