* C:\Users\Bappy\Desktop\Schematic4.sch

* Schematics Version 9.1 - Web Update 1
* Tue Jul 17 09:57:42 2018



** Analysis setup **
.DC LIN V_V1 0V 10V 2 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic4.net"
.INC "Schematic4.als"


.probe


.END
