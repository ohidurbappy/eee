* C:\Users\Bappy\Desktop\PSpiceSchematics\Schematic9.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 25 11:40:46 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic9.net"
.INC "Schematic9.als"


.probe


.END
