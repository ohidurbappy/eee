* C:\Users\Bappy\Desktop\PSpiceSchematics\Schematic7.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 25 11:28:47 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic7.net"
.INC "Schematic7.als"


.probe


.END
