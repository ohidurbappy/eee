* C:\Users\Bappy\Desktop\PSpiceSchematics\Schematic8.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 25 11:37:50 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic8.net"
.INC "Schematic8.als"


.probe


.END
