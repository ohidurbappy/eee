* C:\Users\Bappy\Desktop\Schematic3.sch

* Schematics Version 9.1 - Web Update 1
* Tue Jul 17 09:12:08 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic3.net"
.INC "Schematic3.als"


.probe


.END
