* C:\Users\Bappy\Desktop\PSpiceSchematics\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Sun Nov 25 10:32:33 2018



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
